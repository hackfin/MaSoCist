
module dpram_init_hex_ce_12_32_763e113b4d24162647bd88f925f728963cb7c6a0 #(
	parameter DATA = 32,
	parameter ADDR = 12,
	parameter INIT_HEX = "../sw/bootrom32.hex"
) (

`include "../../common/dpram_hack.vh"

endmodule


